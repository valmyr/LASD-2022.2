module InstrMemory#(parameter WIDTH = 8)(
    input logic  [WIDTH-1:0] address     ,
    output logic [31     :0] RD
);
    
endmodule